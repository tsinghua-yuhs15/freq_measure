module bcd(
  din,
  dout1,
  dout2,
  dout3,
  dout4
);

input   [15:0]   din;
output  [6:0]   dout1,dout2,dout3,dout4;

reg tmp;

assign  dout1=(din[3:0]==4'd0)?7'b1000000:
             (din[3:0]==4'd1)?7'b1111001:
             (din[3:0]==4'd2)?7'b0100100:
             (din[3:0]==4'd3)?7'b0110000:
             (din[3:0]==4'd4)?7'b0011001:
             (din[3:0]==4'd5)?7'b0010010:
             (din[3:0]==4'd6)?7'b0000010:
             (din[3:0]==4'd7)?7'b1111000:
             (din[3:0]==4'd8)?7'b0000000:
             (din[3:0]==4'd9)?7'b0010000:7'b0;

assign  dout2=(din[7:4]==4'd0)?7'b1000000:
             (din[7:4]==4'd1)?7'b1111001:
             (din[7:4]==4'd2)?7'b0100100:
             (din[7:4]==4'd3)?7'b0110000:
             (din[7:4]==4'd4)?7'b0011001:
             (din[7:4]==4'd5)?7'b0010010:
             (din[7:4]==4'd6)?7'b0000010:
             (din[7:4]==4'd7)?7'b1111000:
             (din[7:4]==4'd8)?7'b0000000:
             (din[7:4]==4'd9)?7'b0010000:7'b0;

assign  dout3=(din[11:8]==4'd0)?7'b1000000:
             (din[11:8]==4'd1)?7'b1111001:
             (din[11:8]==4'd2)?7'b0100100:
             (din[11:8]==4'd3)?7'b0110000:
             (din[11:8]==4'd4)?7'b0011001:
             (din[11:8]==4'd5)?7'b0010010:
             (din[11:8]==4'd6)?7'b0000010:
             (din[11:8]==4'd7)?7'b1111000:
             (din[11:8]==4'd8)?7'b0000000:
             (din[11:8]==4'd9)?7'b0010000:7'b0;

assign  dout4=(din[15:12]==4'd0)?7'b1000000:
             (din[15:12]==4'd1)?7'b1111001:
             (din[15:12]==4'd2)?7'b0100100:
             (din[15:12]==4'd3)?7'b0110000:
             (din[15:12]==4'd4)?7'b0011001:
             (din[15:12]==4'd5)?7'b0010010:
             (din[15:12]==4'd6)?7'b0000010:
             (din[15:12]==4'd7)?7'b1111000:
             (din[15:12]==4'd8)?7'b0000000:
             (din[15:12]==4'd9)?7'b0010000:7'b0;
endmodule
